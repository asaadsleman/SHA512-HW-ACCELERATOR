//`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/26/2023 09:51:06 PM
// Design Name: 
// Module Name: k512
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module k512 (
  input [6:0] i,
  output reg [63:0] value
);

  always @*
    case (i)
      0: value = 64'h428a2f98d728ae22;
      1: value = 64'h7137449123ef65cd;
      2: value = 64'hb5c0fbcfec4d3b2f;
      3: value = 64'he9b5dba58189dbbc;
      4: value = 64'h3956c25bf348b538;
      5: value = 64'h59f111f1b605d019;
      6: value = 64'h923f82a4af194f9b;
      7: value = 64'hab1c5ed5da6d8118;
      8: value = 64'hd807aa98a3030242;
      9: value = 64'h12835b0145706fbe;
      10: value = 64'h243185be4ee4b28c;
      11: value = 64'h550c7dc3d5ffb4e2;
      12: value = 64'h72be5d74f27b896f;
      13: value = 64'h80deb1fe3b1696b1;
      14: value = 64'h9bdc06a725c71235;
      15: value = 64'hc19bf174cf692694;
      16: value = 64'he49b69c19ef14ad2;
      17: value = 64'hefbe4786384f25e3;
      18: value = 64'h0fc19dc68b8cd5b5;
      19: value = 64'h240ca1cc77ac9c65;
      20: value = 64'h2de92c6f592b0275;
      21: value = 64'h4a7484aa6ea6e483;
      22: value = 64'h5cb0a9dcbd41fbd4;
      23: value = 64'h76f988da831153b5;
      24: value = 64'h983e5152ee66dfab;
      25: value = 64'ha831c66d2db43210;
      26: value = 64'hb00327c898fb213f;
      27: value = 64'hbf597fc7beef0ee4;
      28: value = 64'hc6e00bf33da88fc2;
      29: value = 64'hd5a79147930aa725;
      30: value = 64'h06ca6351e003826f;
      31: value = 64'h142929670a0e6e70;
      32: value = 64'h27b70a8546d22ffc;
      33: value = 64'h2e1b21385c26c926;
      34: value = 64'h4d2c6dfc5ac42aed;
      35: value = 64'h53380d139d95b3df;
      36: value = 64'h650a73548baf63de;
      37: value = 64'h766a0abb3c77b2a8;
      38: value = 64'h81c2c92e47edaee6;
      39: value = 64'h92722c851482353b;
      40: value = 64'ha2bfe8a14cf10364;
      41: value = 64'ha81a664bbc423001;
      42: value = 64'hc24b8b70d0f89791;
      43: value = 64'hc76c51a30654be30;
      44: value = 64'hd192e819d6ef5218;
      45: value = 64'hd69906245565a910;
      46: value = 64'hf40e35855771202a;
      47: value = 64'h106aa07032bbd1b8;
      48: value = 64'h19a4c116b8d2d0c8;
      49: value = 64'h1e376c085141ab53;
      50: value = 64'h2748774cdf8eeb99;
      51: value = 64'h34b0bcb5e19b48a8;
      52: value = 64'h391c0cb3c5c95a63;
      53: value = 64'h4ed8aa4ae3418acb;
      54: value = 64'h5b9cca4f7763e373;
      55: value = 64'h682e6ff3d6b2b8a3;
      56: value = 64'h748f82ee5defb2fc;
      57: value = 64'h78a5636f43172f60;
      58: value = 64'h84c87814a1f0ab72;
      59: value = 64'h8cc702081a6439ec;
      60: value = 64'h90befffa23631e28;
      61: value = 64'ha4506cebde82bde9;
      62: value = 64'hbef9a3f7b2c67915;
      63: value = 64'hc67178f2e372532b;
      64: value = 64'hca273eceea26619c;
      65: value = 64'hd186b8c721c0c207;
      66: value = 64'heada7dd6cde0eb1e;
      67: value = 64'hf57d4f7fee6ed178;
      68: value = 64'h06f067aa72176fba;
      69: value = 64'h0a637dc5a2c898a6;
      70: value = 64'h113f9804bef90dae;
      71: value = 64'h1b710b35131c471b;
      72: value = 64'h28db77f523047d84;
      73: value = 64'h32caab7b40c72493;
      74: value = 64'h3c9ebe0a15c9bebc;
      75: value = 64'h431d67c49c100d4c;
      76: value = 64'h4cc5d4becb3e42b6;
      77: value = 64'h597f299cfc657e2a;
      78: value = 64'h5fcb6fab3ad6faec;
      79: value = 64'h6c44198c4a475817;
      default: value = 64'h0;
    endcase

endmodule

